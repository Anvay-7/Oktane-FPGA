module fpga (
	inout  [23:0] p    ,
	input         sin  ,
	input         s_clk,
	input         f_clk,
	input         flag ,
	output        sout
);
	wire v000,v001,v002,v003;
	wire v010,v011,v012,v013;
	wire v020,v021,v022,v023;
	wire v030,v031,v032,v033;
	wire v100,v101,v102,v103;
	wire v110,v111,v112,v113;
	wire v120,v121,v122,v123;
	wire v130,v131,v132,v133;
	wire v200,v201,v202,v203;
	wire v210,v211,v212,v213;
	wire v220,v221,v222,v223;
	wire v230,v231,v232,v233;

	wire h000,h001,h002,h003;
	wire h010,h011,h012,h013;
	wire h020,h021,h022,h023;
	wire h100,h101,h102,h103;
	wire h110,h111,h112,h113;
	wire h120,h121,h122,h123;
	wire h200,h201,h202,h203;
	wire h210,h211,h212,h213;
	wire h220,h221,h222,h223;
	wire h300,h301,h302,h303;
	wire h310,h311,h312,h313;
	wire h320,h321,h322,h323;

	wire y01, y02, y11, y12, y21, y22, y31, y32, y41, y42, y51, y52, y61, y62, y71, y72, y81, y82;

	assign sys_clk = s_clk & flag;
	
	assign y01 = (!flag) ? y01_clb : 1'bz;
	assign y02 = (!flag) ? y02_clb : 1'bz;
	assign y11 = (!flag) ? y11_clb : 1'bz;
	assign y12 = (!flag) ? y12_clb : 1'bz;
	assign y21 = (!flag) ? y21_clb : 1'bz;
	assign y22 = (!flag) ? y22_clb : 1'bz;
	assign y31 = (!flag) ? y31_clb : 1'bz;
	assign y32 = (!flag) ? y32_clb : 1'bz;
	assign y41 = (!flag) ? y41_clb : 1'bz;
	assign y42 = (!flag) ? y42_clb : 1'bz;
	assign y51 = (!flag) ? y51_clb : 1'bz;
	assign y52 = (!flag) ? y52_clb : 1'bz;
	assign y61 = (!flag) ? y61_clb : 1'bz;
	assign y62 = (!flag) ? y62_clb : 1'bz;
	assign y71 = (!flag) ? y71_clb : 1'bz;
	assign y72 = (!flag) ? y72_clb : 1'bz;
	assign y81 = (!flag) ? y81_clb : 1'bz;
	assign y82 = (!flag) ? y82_clb : 1'bz;


	switch_box s_00 (.l(), .u(), .r(h000), .d(v000), .clk(sys_clk), .si(sin), .so(s01));
	switch_box s_01 (.l(), .u(), .r(h001), .d(v001), .clk(sys_clk), .si(s01), .so(s02));
	switch_box s_02 (.l(), .u(), .r(h002), .d(v002), .clk(sys_clk), .si(s02), .so(s03));
	switch_box s_03 (.l(), .u(), .r(h003), .d(v003), .clk(sys_clk), .si(s03), .so(c23));

	/////////////////////////////////////////////////////////////////////////////////////////
	conn_box c_23 (.a({h003,h002,h001,h000}), .b(p[23]), .clk(sys_clk), .si(c23), .so(c22));
	conn_box c_22 (.a({h003,h002,h001,h000}), .b(p[22]), .clk(sys_clk), .si(c22), .so(s10));

	/////////////////////////////////////////////////////////////////////////////////////////
	switch_box s_10 (.l(h000), .u(), .r(h010), .d(v010), .clk(sys_clk), .si(s10), .so(s11));
	switch_box s_11 (.l(h001), .u(), .r(h011), .d(v011), .clk(sys_clk), .si(s11), .so(s12));
	switch_box s_12 (.l(h002), .u(), .r(h012), .d(v012), .clk(sys_clk), .si(s12), .so(s13));
	switch_box s_13 (.l(h003), .u(), .r(h013), .d(v013), .clk(sys_clk), .si(s13), .so(c21));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_21 (.a({h013,h012,h011,h010}), .b(p[21]), .clk(sys_clk), .si(c21), .so(c20));
	conn_box c_20 (.a({h013,h012,h011,h010}), .b(p[20]), .clk(sys_clk), .si(c20), .so(s20));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_20 (.l(h010), .u(), .r(h020), .d(v020), .clk(sys_clk), .si(s20), .so(s21));
	switch_box s_21 (.l(h011), .u(), .r(h021), .d(v021), .clk(sys_clk), .si(s21), .so(s22));
	switch_box s_22 (.l(h012), .u(), .r(h022), .d(v022), .clk(sys_clk), .si(s22), .so(s23));
	switch_box s_23 (.l(h013), .u(), .r(h023), .d(v023), .clk(sys_clk), .si(s23), .so(c19));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_19 (.a({h023,h022,h021,h020}), .b(p[19]), .clk(sys_clk), .si(c19), .so(c18));
	conn_box c_18 (.a({h023,h022,h021,h020}), .b(p[18]), .clk(sys_clk), .si(c18), .so(s30));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_30 (.l(h020), .u(), .r(h030), .d(v030), .clk(sys_clk), .si(s30), .so(s31));
	switch_box s_31 (.l(h021), .u(), .r(h031), .d(v031), .clk(sys_clk), .si(s31), .so(s32));
	switch_box s_32 (.l(h022), .u(), .r(h032), .d(v032), .clk(sys_clk), .si(s32), .so(s33));
	switch_box s_33 (.l(h023), .u(), .r(h033), .d(v033), .clk(sys_clk), .si(s33), .so(c28));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_28 (.a({v030,v031,v032,v033}), .b(y21), .clk(sys_clk), .si(c28), .so(c17));

	conn_box c_17 (.a({v033,v032,v031,v030}), .b(p[17]), .clk(sys_clk), .si(c17), .so(c16));
	conn_box c_16 (.a({v033,v032,v031,v030}), .b(p[16]), .clk(sys_clk), .si(c16), .so(c29));

	conn_box c_29 (.a({v030,v031,v032,v033}), .b(y22), .clk(sys_clk), .si(c29), .so(d2));

	/////////////////////////////////////////////////////////////////////////////////////////

	clb slice_2 (.si(d2), .sys_clk(sys_clk), .a({v023,v022,v021,v020}), .b({h023,h022,h021,h020}), .c({h123,h122,h121,h120}), .clk({h122,h121,h120}), .f_clk(f_clk), .y1(y21_clb), .y2(y22_clb), .so(c26));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_26 (.a({v020,v021,v022,v023}), .b(y11), .clk(sys_clk), .si(c26), .so(c27));
	conn_box c_27 (.a({v020,v021,v022,v023}), .b(y12), .clk(sys_clk), .si(c27), .so(d1));

	/////////////////////////////////////////////////////////////////////////////////////////

	clb slice_1 (.si(d1), .sys_clk(sys_clk), .a({v013,v012,v011,v010}), .b({h013,h012,h011,h010}), .c({h113,h112,h111,h110}), .clk({h112,h111,h110}), .f_clk(f_clk), .y1(y11_clb), .y2(y12_clb), .so(c24));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_24 (.a({v010,v011,v012,v013}), .b(y01), .clk(sys_clk), .si(c24), .so(c25));
	conn_box c_25 (.a({v010,v011,v012,v013}), .b(y02), .clk(sys_clk), .si(c25), .so(d0));

	/////////////////////////////////////////////////////////////////////////////////////////

	clb slice_0 (.si(d0), .sys_clk(sys_clk), .a({v003,v002,v001,v000}), .b({h003,h002,h001,h000}), .c({h103,h102,h101,h100}), .clk({h102,h101,h100}), .f_clk(f_clk), .y1(y01_clb), .y2(y02_clb), .so(c0));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_0 (.a({v000,v001,v002,v003}), .b(p[0]), .clk(sys_clk), .si(c0), .so(c1));
	conn_box c_1 (.a({v000,v001,v002,v003}), .b(p[1]), .clk(sys_clk), .si(c1), .so(s40));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_40 (.l(), .u(v000), .r(h100), .d(v100), .clk(sys_clk), .si(s40), .so(s41));
	switch_box s_41 (.l(), .u(v001), .r(h101), .d(v101), .clk(sys_clk), .si(s41), .so(s42));
	switch_box s_42 (.l(), .u(v002), .r(h102), .d(v102), .clk(sys_clk), .si(s42), .so(s43));
	switch_box s_43 (.l(), .u(v003), .r(h103), .d(v103), .clk(sys_clk), .si(s43), .so(s50));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_50 (.l(h100), .u(v010), .r(h110), .d(v110), .clk(sys_clk), .si(s50), .so(s51));
	switch_box s_51 (.l(h101), .u(v011), .r(h111), .d(v111), .clk(sys_clk), .si(s51), .so(s52));
	switch_box s_52 (.l(h102), .u(v012), .r(h112), .d(v112), .clk(sys_clk), .si(s52), .so(s53));
	switch_box s_53 (.l(h103), .u(v013), .r(h113), .d(v113), .clk(sys_clk), .si(s53), .so(s60));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_60 (.l(h110), .u(v020), .r(h120), .d(v120), .clk(sys_clk), .si(s60), .so(s61));
	switch_box s_61 (.l(h111), .u(v021), .r(h121), .d(v121), .clk(sys_clk), .si(s61), .so(s62));
	switch_box s_62 (.l(h112), .u(v022), .r(h122), .d(v122), .clk(sys_clk), .si(s62), .so(s63));
	switch_box s_63 (.l(h113), .u(v023), .r(h123), .d(v123), .clk(sys_clk), .si(s63), .so(s70));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_70 (.l(h120), .u(v030), .r(), .d(v130), .clk(sys_clk), .si(s70), .so(s71));
	switch_box s_71 (.l(h121), .u(v031), .r(), .d(v131), .clk(sys_clk), .si(s71), .so(s72));
	switch_box s_72 (.l(h122), .u(v032), .r(), .d(v132), .clk(sys_clk), .si(s72), .so(s73));
	switch_box s_73 (.l(h123), .u(v033), .r(), .d(v133), .clk(sys_clk), .si(s73), .so(c34));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_34 (.a({v130,v131,v132,v133}), .b(y51), .clk(sys_clk), .si(c34), .so(c15));

	conn_box c_15 (.a({v130,v131,v132,v133}), .b(p[15]), .clk(sys_clk), .si(c15), .so(c14));
	conn_box c_14 (.a({v130,v131,v132,v133}), .b(p[14]), .clk(sys_clk), .si(c14), .so(c35));

	conn_box c_35 (.a({v130,v131,v132,v133}), .b(y52), .clk(sys_clk), .si(c35), .so(d5));

	/////////////////////////////////////////////////////////////////////////////////////////

	clb slice_5 (.si(d5), .sys_clk(sys_clk), .a({v123,v122,v121,v120}), .b({h123,h122,h121,h120}), .c({h223,h222,h221,h220}), .clk({h222,h221,h220}), .f_clk(f_clk), .y1(y51_clb), .y2(y52_clb), .so(c32));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_32 (.a({v120,v121,v122,v123}), .b(y41), .clk(sys_clk), .si(c32), .so(c33));
	conn_box c_33 (.a({v120,v121,v122,v123}), .b(y42), .clk(sys_clk), .si(c33), .so(d4));

	/////////////////////////////////////////////////////////////////////////////////////////

	clb slice_4 (.si(d4), .sys_clk(sys_clk), .a({v113,v112,v111,v110}), .b({h113,h112,h111,h110}), .c({h213,h212,h211,h210}), .clk({h212,h211,h210}), .f_clk(f_clk), .y1(y41_clb), .y2(y42_clb), .so(c30));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_30 (.a({v110,v111,v112,v113}), .b(y31), .clk(sys_clk), .si(c30), .so(c31));
	conn_box c_31 (.a({v110,v111,v112,v113}), .b(y32), .clk(sys_clk), .si(c31), .so(d3));

	/////////////////////////////////////////////////////////////////////////////////////////

	clb slice_3 (.si(d3), .sys_clk(sys_clk), .a({v103,v102,v101,v100}), .b({h103,h102,h101,h100}), .c({h203,h202,h201,h200}), .clk({h202,h201,h200}), .f_clk(f_clk), .y1(y31_clb), .y2(y32_clb), .so(c2));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_2 (.a({v100,v101,v102,v103}), .b(p[2]), .clk(sys_clk), .si(c2), .so(c3));
	conn_box c_3 (.a({v100,v101,v102,v103}), .b(p[3]), .clk(sys_clk), .si(c3), .so(s80));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_80 (.l(), .u(v100), .r(h200), .d(v200), .clk(sys_clk), .si(s80), .so(s81));
	switch_box s_81 (.l(), .u(v101), .r(h201), .d(v201), .clk(sys_clk), .si(s81), .so(s82));
	switch_box s_82 (.l(), .u(v102), .r(h202), .d(v202), .clk(sys_clk), .si(s82), .so(s83));
	switch_box s_83 (.l(), .u(v103), .r(h203), .d(v203), .clk(sys_clk), .si(s83), .so(s90));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_90 (.l(h200), .u(v110), .r(h210), .d(v210), .clk(sys_clk), .si(s90), .so(s91));
	switch_box s_91 (.l(h201), .u(v111), .r(h211), .d(v211), .clk(sys_clk), .si(s91), .so(s92));
	switch_box s_92 (.l(h202), .u(v112), .r(h212), .d(v212), .clk(sys_clk), .si(s92), .so(s93));
	switch_box s_93 (.l(h203), .u(v113), .r(h213), .d(v213), .clk(sys_clk), .si(s93), .so(s100));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_100 (.l(h210), .u(v120), .r(h220), .d(v220), .clk(sys_clk), .si(s100), .so(s101));
	switch_box s_101 (.l(h211), .u(v121), .r(h221), .d(v221), .clk(sys_clk), .si(s101), .so(s102));
	switch_box s_102 (.l(h212), .u(v122), .r(h222), .d(v222), .clk(sys_clk), .si(s102), .so(s103));
	switch_box s_103 (.l(h213), .u(v123), .r(h223), .d(v223), .clk(sys_clk), .si(s103), .so(s110));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_110 (.l(h220), .u(v130), .r(), .d(v230), .clk(sys_clk), .si(s110), .so(s111));
	switch_box s_111 (.l(h221), .u(v131), .r(), .d(v231), .clk(sys_clk), .si(s111), .so(s112));
	switch_box s_112 (.l(h222), .u(v132), .r(), .d(v232), .clk(sys_clk), .si(s112), .so(s113));
	switch_box s_113 (.l(h223), .u(v133), .r(), .d(v233), .clk(sys_clk), .si(s113), .so(c40));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_40 (.a({v230,v231,v232,v233}), .b(y81), .clk(sys_clk), .si(c40), .so(c13));

	conn_box c_13 (.a({v230,v231,v232,v233}), .b(p[13]), .clk(sys_clk), .si(c13), .so(c12));
	conn_box c_12 (.a({v230,v231,v232,v233}), .b(p[12]), .clk(sys_clk), .si(c12), .so(c41));

	conn_box c_41 (.a({v230,v231,v232,v233}), .b(y82), .clk(sys_clk), .si(c41), .so(d8));

	/////////////////////////////////////////////////////////////////////////////////////////

	clb slice_8 (.si(d8), .sys_clk(sys_clk), .a({v223,v222,v221,v220}), .b({h223,h222,h221,h220}), .c({h323,h322,h321,h320}), .clk({h322,h321,h320}), .f_clk(f_clk), .y1(y81_clb), .y2(y82_clb), .so(c38));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_38 (.a({v220,v221,v222,v223}), .b(y71), .clk(sys_clk), .si(c38), .so(c39));
	conn_box c_39 (.a({v220,v221,v222,v223}), .b(y72), .clk(sys_clk), .si(c39), .so(d7));

	/////////////////////////////////////////////////////////////////////////////////////////

	clb slice_7 (.si(d7), .sys_clk(sys_clk), .a({v213,v212,v211,v210}), .b({h213,h212,h211,h210}), .c({h313,h312,h311,h310}), .clk({h312,h311,h310}), .f_clk(f_clk), .y1(y71_clb), .y2(y72_clb), .so(c36));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_36 (.a({v210,v211,v212,v213}), .b(y61), .clk(sys_clk), .si(c36), .so(c37));
	conn_box c_37 (.a({v210,v211,v212,v213}), .b(y62), .clk(sys_clk), .si(c37), .so(d6));

	/////////////////////////////////////////////////////////////////////////////////////////

	clb slice_6 (.si(d6), .sys_clk(sys_clk), .a({v203,v202,v201,v200}), .b({h203,h202,h201,h200}), .c({h303,h302,h301,h300}), .clk({h302,h301,h300}), .f_clk(f_clk), .y1(y61_clb), .y2(y62_clb), .so(c4));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_4 (.a({v200,v201,v202,v203}), .b(p[4]), .clk(sys_clk), .si(c4), .so(c5));
	conn_box c_5 (.a({v200,v201,v202,v203}), .b(p[5]), .clk(sys_clk), .si(c5), .so(s120));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_120 (.l(), .u(v200), .r(h300), .d(), .clk(sys_clk), .si(s120), .so(s121));
	switch_box s_121 (.l(), .u(v201), .r(h301), .d(), .clk(sys_clk), .si(s121), .so(s122));
	switch_box s_122 (.l(), .u(v202), .r(h302), .d(), .clk(sys_clk), .si(s122), .so(s123));
	switch_box s_123 (.l(), .u(v203), .r(h303), .d(), .clk(sys_clk), .si(s123), .so(c6));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_6 (.a({h300,h301,h302,h303}), .b(p[6]), .clk(sys_clk), .si(c6), .so(c7));
	conn_box c_7 (.a({h300,h301,h302,h303}), .b(p[7]), .clk(sys_clk), .si(c7), .so(s130));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_130 (.l(h300), .u(v210), .r(h310), .d(), .clk(sys_clk), .si(s130), .so(s131));
	switch_box s_131 (.l(h301), .u(v211), .r(h311), .d(), .clk(sys_clk), .si(s131), .so(s132));
	switch_box s_132 (.l(h302), .u(v212), .r(h312), .d(), .clk(sys_clk), .si(s132), .so(s133));
	switch_box s_133 (.l(h303), .u(v213), .r(h313), .d(), .clk(sys_clk), .si(s133), .so(c8));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_8 (.a({h310,h311,h312,h313}), .b(p[8]), .clk(sys_clk), .si(c8), .so(c9));
	conn_box c_9 (.a({h310,h311,h312,h313}), .b(p[9]), .clk(sys_clk), .si(c9), .so(s140));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_140 (.l(h310), .u(v220), .r(h320), .d(), .clk(sys_clk), .si(s140), .so(s141));
	switch_box s_141 (.l(h311), .u(v221), .r(h321), .d(), .clk(sys_clk), .si(s141), .so(s142));
	switch_box s_142 (.l(h312), .u(v222), .r(h322), .d(), .clk(sys_clk), .si(s142), .so(s143));
	switch_box s_143 (.l(h313), .u(v223), .r(h323), .d(), .clk(sys_clk), .si(s143), .so(c10));

	/////////////////////////////////////////////////////////////////////////////////////////

	conn_box c_10 (.a({h320,h321,h322,h323}), .b(p[10]), .clk(sys_clk), .si(c10), .so(c11));
	conn_box c_11 (.a({h320,h321,h322,h323}), .b(p[11]), .clk(sys_clk), .si(c11), .so(s150));

	/////////////////////////////////////////////////////////////////////////////////////////

	switch_box s_150 (.l(h320), .u(v230), .r(), .d(), .clk(sys_clk), .si(s150), .so(s151));
	switch_box s_151 (.l(h321), .u(v231), .r(), .d(), .clk(sys_clk), .si(s151), .so(s152));
	switch_box s_152 (.l(h322), .u(v232), .r(), .d(), .clk(sys_clk), .si(s152), .so(s153));
	switch_box s_153 (.l(h323), .u(v233), .r(), .d(), .clk(sys_clk), .si(s153), .so(sout));

endmodule
